module cpu();



endmodule
